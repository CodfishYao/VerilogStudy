module adder_tb();
endmodule