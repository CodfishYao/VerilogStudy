module mul_tc_16_16(
    input [15:0] a,
    input [15:0] b,
    output[31:0] product
);

endmodule